interface operation;
  logic d,clk,rst;
  logic q,qb;
 endinterface
