class transaction;
  rand logic d;
   logic clk;
  //logic d;
   logic rst;
  bit q;
  bit qb;
endclass
